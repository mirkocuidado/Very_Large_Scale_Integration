library verilog;
use verilog.vl_types.all;
entity top_t_ff is
end top_t_ff;
