library verilog;
use verilog.vl_types.all;
entity lab1_kombinaciona_testbench is
end lab1_kombinaciona_testbench;
