library verilog;
use verilog.vl_types.all;
entity top_register is
end top_register;
