library verilog;
use verilog.vl_types.all;
entity lab1_sekvencijalna_testbench is
end lab1_sekvencijalna_testbench;
