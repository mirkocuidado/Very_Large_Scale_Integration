library verilog;
use verilog.vl_types.all;
entity dut is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        \in\            : in     vl_logic_vector(3 downto 0);
        ctrl            : in     vl_logic_vector(2 downto 0);
        \out\           : out    vl_logic_vector(3 downto 0)
    );
end dut;
