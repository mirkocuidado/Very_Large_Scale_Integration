library verilog;
use verilog.vl_types.all;
entity top_jk_ff is
end top_jk_ff;
