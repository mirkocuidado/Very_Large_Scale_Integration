library verilog;
use verilog.vl_types.all;
entity top_d_ff is
end top_d_ff;
